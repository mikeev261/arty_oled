`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03/03/2017 10:44:57 PM
// Design Name: 
// Module Name: oled_ctrl
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments: https://reference.digilentinc.com/_media/reference/pmod/pmodoledrgb/pmodoledrgb_rm.pdf
// 
//////////////////////////////////////////////////////////////////////////////////


module oled_ctrl(

    );
endmodule